library ieee;
use ieee.std_logic_1164.all;
entity song is
port
(
	clk8hz						:in std_logic;--12MHz
	tone2						:out integer range 0 to 10;
	music_num					:in std_logic;
	num    						:in integer range 0 to 1
);
end entity;

architecture song_arch of song is
signal ptr    :integer range 0 to 228;
begin
process(clk8hz, music_num, num)
begin
if music_num='1' then ptr <= 0;  --After pushing the button, switch tune immediately.
else
if rising_edge(clk8hz) then--ÿ0.125s�任����
  if ptr = 228 then ptr <= 0;
  else ptr <= ptr + 1;
  end if;
case num is
when 0=>                         --Music No.1 Twinkle Twinkle Little Star
  case ptr is
when	1	=>tone2 <=	1	;--do
when	2	=>tone2 <=	1	;
when	3	=>tone2 <=	1	;
when	4	=>tone2 <=	1	;
when	5	=>tone2 <=	0	;
when	6	=>tone2 <=	1	;
when	7	=>tone2 <=	1	;
when	8	=>tone2 <=	1	;
when	9	=>tone2 <=	1	;
when	10	=>tone2 <=	0	;
when	11	=>tone2 <=	5	;
when	12	=>tone2 <=	5	;
when	13	=>tone2 <=	5	;
when	14	=>tone2 <=	5	;
when	15	=>tone2 <=	0	;
when	16	=>tone2 <=	5	;
when	17	=>tone2 <=	5	;
when	18	=>tone2 <=	5	;
when	19	=>tone2 <=	5	;
when	20	=>tone2 <=	0	;
when	21	=>tone2 <=	6	;
when	22	=>tone2 <=	6	;
when	23	=>tone2 <=	6	;
when	24	=>tone2 <=	6	;
when	25	=>tone2 <=	0	;
when	26	=>tone2 <=	6	;
when	27	=>tone2 <=	6	;
when	28	=>tone2 <=	6	;
when	29	=>tone2 <=	6	;
when	30	=>tone2 <=	0	;
when	31	=>tone2 <=	5	;
when	32	=>tone2 <=	5	;
when	33	=>tone2 <=	5	;
when	34	=>tone2 <=	5	;
when	35	=>tone2 <=	0	;
when	36	=>tone2 <=	0	;
when	37	=>tone2 <=	0	;
when	38	=>tone2<=	0	;
when	39	=>tone2<=	4	;
when	40	=>tone2<=	4	;
when	41	=>tone2<=	4	;
when	42	=>tone2<=	4	;
when	43	=>tone2<=	0	;
when	44	=>tone2<=	4	;
when	45	=>tone2<=	4	;
when	46	=>tone2<=	4	;
when	47	=>tone2<=	4	;
when	48	=>tone2<=	0	;
when	49	=>tone2<=	3	;
when	50	=>tone2<=	3	;
when	51	=>tone2<=	3	;
when	52	=>tone2<=	3	;
when	53	=>tone2<=	0	;
when	54	=>tone2<=	3	;
when	55	=>tone2<=	3	;
when	56	=>tone2<=	3	;
when	57	=>tone2<=	3	;
when	58	=>tone2<=	0	;
when	59	=>tone2<=	2	;
when	60	=>tone2<=	2	;
when	61	=>tone2<=	2	;
when	62	=>tone2<=	2	;
when	63	=>tone2<=	0	;
when	64	=>tone2<=	2	;
when	65	=>tone2<=	2	;
when	66	=>tone2<=	2	;
when	67	=>tone2<=	2	;
when	68	=>tone2<=	0	;
when	69	=>tone2<=	1	;
when	70	=>tone2<=	1	;
when	71	=>tone2<=	1	;
when	72	=>tone2<=	1	;
when	73	=>tone2<=	0	;
when	74	=>tone2<=	0	;
when	75	=>tone2<=	0	;
when	76	=>tone2<=	0	;
when	77	=>tone2<=	5	;
when	78	=>tone2<=	5	;
when	79	=>tone2<=	5	;
when	80	=>tone2<=	5	;
when	81	=>tone2<=	0	;
when	82	=>tone2<=	5	;
when	83	=>tone2<=	5	;
when	84	=>tone2<=	5	;
when	85	=>tone2<=	5	;
when	86	=>tone2<=	0	;
when	87	=>tone2<=	4	;
when	88	=>tone2<=	4	;
when	89	=>tone2<=	4	;
when	90	=>tone2<=	4	;
when	91	=>tone2<=	0	;
when	92	=>tone2<=	4	;
when	93	=>tone2<=	4	;
when	94	=>tone2<=	4	;
when	95	=>tone2<=	4	;
when	96	=>tone2<=	0	;
when	97	=>tone2<=	3	;
when	98	=>tone2<=	3	;
when	99	=>tone2<=	3	;
when	100	=>tone2<=	3	;
when	101	=>tone2<=	0	;
when	102	=>tone2<=	3	;
when	103	=>tone2<=	3	;
when	104	=>tone2<=	3	;
when	105	=>tone2<=	3	;
when	106	=>tone2<=	0	;
when	107	=>tone2<=	2	;
when	108	=>tone2<=	2	;
when	109	=>tone2<=	2	;
when	110	=>tone2<=	2	;
when	111	=>tone2<=	0	;
when	112	=>tone2<=	0	;
when	113	=>tone2<=	0	;
when	114	=>tone2<=	0	;
when	115	=>tone2<=	5	;
when	116	=>tone2<=	5	;
when	117	=>tone2<=	5	;
when	118	=>tone2<=	5	;
when	119	=>tone2<=	0	;
when	120	=>tone2<=	5	;
when	121	=>tone2<=	5	;
when	122	=>tone2<=	5	;
when	123	=>tone2<=	5	;
when	124	=>tone2<=	0	;
when	125	=>tone2<=	4	;
when	126	=>tone2<=	4	;
when	127	=>tone2<=	4	;
when	128	=>tone2<=	4	;
when	129	=>tone2<=	0	;
when	130	=>tone2<=	4	;
when	131	=>tone2<=	4	;
when	132	=>tone2<=	4	;
when	133	=>tone2<=	4	;
when	134	=>tone2<=	0	;
when	135	=>tone2<=	3	;
when	136	=>tone2<=	3	;
when	137	=>tone2<=	3	;
when	138	=>tone2<=	3	;
when	139	=>tone2<=	0	;
when	140	=>tone2<=	3	;
when	141	=>tone2<=	3	;
when	142	=>tone2<=	3	;
when	143	=>tone2<=	3	;
when	144	=>tone2<=	0	;
when	145	=>tone2<=	2	;
when	146	=>tone2<=	2	;
when	147	=>tone2<=	2	;
when	148	=>tone2<=	2	;
when	149	=>tone2<=	0	;
when	150	=>tone2<=	0	;
when	151	=>tone2<=	0	;
when	152	=>tone2<=	0	;
when	153	=>tone2<=	1	;
when	154	=>tone2<=	1	;
when	155	=>tone2<=	1	;
when	156	=>tone2<=	1	;
when	157	=>tone2<=	0	;
when	158	=>tone2<=	1	;
when	159	=>tone2<=	1	;
when	160	=>tone2<=	1	;
when	161	=>tone2<=	1	;
when	162	=>tone2<=	0	;
when	163	=>tone2<=	5	;
when	164	=>tone2<=	5	;
when	165	=>tone2<=	5	;
when	166	=>tone2<=	5	;
when	167	=>tone2<=	0	;
when	168	=>tone2<=	5	;
when	169	=>tone2<=	5	;
when	170	=>tone2<=	5	;
when	171	=>tone2<=	5	;
when	172	=>tone2<=	0	;
when	173	=>tone2<=	6	;
when	174	=>tone2<=	6	;
when	175	=>tone2<=	6	;
when	176	=>tone2<=	6	;
when	177	=>tone2<=	0	;
when	178	=>tone2<=	6	;
when	179	=>tone2<=	6	;
when	180	=>tone2<=	6	;
when	181	=>tone2<=	6	;
when	182	=>tone2<=	0	;
when	183	=>tone2<=	5	;
when	184	=>tone2<=	5	;
when	185	=>tone2<=	5	;
when	186	=>tone2<=	5	;
when	187	=>tone2<=	0	;
when	188	=>tone2<=	0	;
when	189	=>tone2<=	0	;
when	190	=>tone2<=	0	;
when	191	=>tone2<=	4	;
when	192	=>tone2<=	4	;
when	193	=>tone2<=	4	;
when	194	=>tone2<=	4	;
when	195	=>tone2<=	0	;
when	196	=>tone2<=	4	;
when	197	=>tone2<=	4	;
when	198	=>tone2<=	4	;
when	199	=>tone2<=	4	;
when	200	=>tone2<=	0	;
when	201	=>tone2<=	3	;
when	202	=>tone2<=	3	;
when	203	=>tone2<=	3	;
when	204	=>tone2<=	3	;
when	205	=>tone2<=	0	;
when	206	=>tone2<=	3	;
when	207	=>tone2<=	3	;
when	208	=>tone2<=	3	;
when	209	=>tone2<=	3	;
when	210	=>tone2<=	0	;
when	211	=>tone2<=	2	;
when	212	=>tone2<=	2	;
when	213	=>tone2<=	2	;
when	214	=>tone2<=	2	;
when	215	=>tone2<=	0	;
when	216	=>tone2<=	2	;
when	217	=>tone2<=	2	;
when	218	=>tone2<=	2	;
when	219	=>tone2<=	2	;
when	220	=>tone2<=	0	;
when	221	=>tone2<=	1	;
when	222	=>tone2<=	1	;
when	223	=>tone2<=	1	;
when	224	=>tone2<=	1	;
when	225	=>tone2<=	0	;
when	226	=>tone2<=	0	;
when	227	=>tone2<=	0	;
when	228	=>tone2<=	0	;
  when others =>tone2<=0;
  end case;
when 1=>                --Music 2
 case ptr is
when	1	=>tone2<=	6	;
when	2	=>tone2<=	6	;
when	3	=>tone2<=	0	;
when	4	=>tone2<=	7	;
when	5	=>tone2<=	7	;
when	6	=>tone2<=	0	;
when	7	=>tone2<=	8	;
when	8	=>tone2<=	8	;
when	9	=>tone2<=	8	;
when	10	=>tone2<=	8	;
when	11	=>tone2<=	0	;
when	12	=>tone2<=	7	;
when	13	=>tone2<=	7	;
when	14	=>tone2<=	0	;
when	15	=>tone2<=	8	;
when	16	=>tone2<=	8	;
when	17	=>tone2<=	8	;
when	18	=>tone2<=	8	;
when	19	=>tone2<=	0	;
when	20	=>tone2<=	10	;
when	21	=>tone2<=	10	;
when	22	=>tone2<=	10	;
when	23	=>tone2<=	10	;
when	24	=>tone2<=	0	;
when	25	=>tone2<=	7	;
when	26	=>tone2<=	7	;
when	27	=>tone2<=	7	;
when	28	=>tone2<=	7	;
when	29	=>tone2<=	7	;
when	30	=>tone2<=	7	;
when	31	=>tone2<=	0	;
when	32	=>tone2<=	3	;
when	33	=>tone2<=	3	;
when	34	=>tone2<=	3	;
when	35	=>tone2<=	3	;
when	36	=>tone2<=	0	;
when	37	=>tone2<=	6	;
when	38	=>tone2<=	6	;
when	39	=>tone2<=	6	;
when	40	=>tone2<=	6	;
when	41	=>tone2<=	6	;
when	42	=>tone2<=	6	;
when	43	=>tone2<=	0	;
when	44	=>tone2<=	5	;
when	45	=>tone2<=	5	;
when	46	=>tone2<=	0	;
when	47	=>tone2<=	6	;
when	48	=>tone2<=	6	;
when	49	=>tone2<=	6	;
when	50	=>tone2<=	6	;
when	51	=>tone2<=	0	;
when	52	=>tone2<=	8	;
when	53	=>tone2<=	8	;
when	54	=>tone2<=	8	;
when	55	=>tone2<=	8	;
when	56	=>tone2<=	0	;
when	57	=>tone2<=	5	;
when	58	=>tone2<=	5	;
when	59	=>tone2<=	5	;
when	60	=>tone2<=	5	;
when	61	=>tone2<=	5	;
when	62	=>tone2<=	5	;
when	63	=>tone2<=	0	;
when	64	=>tone2<=	2	;
when	65	=>tone2<=	2	;
when	66	=>tone2<=	0	;
when	67	=>tone2<=	3	;
when	68	=>tone2<=	3	;
when	69	=>tone2<=	0	;
when	70	=>tone2<=	4	;
when	71	=>tone2<=	4	;
when	72	=>tone2<=	4	;
when	73	=>tone2<=	4	;
when	74	=>tone2<=	4	;
when	75	=>tone2<=	4	;
when	76	=>tone2<=	0	;
when	77	=>tone2<=	3	;
when	78	=>tone2<=	3	;
when	79	=>tone2<=	0	;
when	80	=>tone2<=	4	;
when	81	=>tone2<=	4	;
when	82	=>tone2<=	0	;
when	83	=>tone2<=	8	;
when	84	=>tone2<=	8	;
when	85	=>tone2<=	8	;
when	86	=>tone2<=	8	;
when	87	=>tone2<=	8	;
when	88	=>tone2<=	8	;
when	89	=>tone2<=	0	;
when	90	=>tone2<=	3	;
when	91	=>tone2<=	3	;
when	92	=>tone2<=	3	;
when	93	=>tone2<=	3	;
when	94	=>tone2<=	3	;
when	95	=>tone2<=	3	;
when	96	=>tone2<=	0	;
when	97	=>tone2<=	2	;
when	98	=>tone2<=	2	;
when	99	=>tone2<=	0	;
when	100	=>tone2<=	3	;
when	101	=>tone2<=	3	;
when	102	=>tone2<=	0	;
when	103	=>tone2<=	8	;
when	104	=>tone2<=	8	;
when	105	=>tone2<=	8	;
when	106	=>tone2<=	8	;
when	107	=>tone2<=	8	;
when	108	=>tone2<=	8	;
when	109	=>tone2<=	0	;
when	110	=>tone2<=	7	;
when	111	=>tone2<=	7	;
when	112	=>tone2<=	7	;
when	113	=>tone2<=	7	;
when	114	=>tone2<=	7	;
when	115	=>tone2<=	0	;
when	116	=>tone2<=	5	;
when	117	=>tone2<=	5	;
when	118	=>tone2<=	0	;
when	119	=>tone2<=	5	;
when	120	=>tone2<=	5	;
when	121	=>tone2<=	5	;
when	122	=>tone2<=	0	;
when	123	=>tone2<=	7	;
when	124	=>tone2<=	7	;
when	125	=>tone2<=	7	;
when	126	=>tone2<=	7	;
when	127	=>tone2<=	0	;
when	128	=>tone2<=	7	;
when	129	=>tone2<=	7	;
when	130	=>tone2<=	7	;
when	131	=>tone2<=	7	;
when	132	=>tone2<=	7	;
when	133	=>tone2<=	7	;
when	134	=>tone2<=	0	;
when	135	=>tone2<=	6	;
when	136	=>tone2<=	6	;
when	137	=>tone2<=	0	;
when	138	=>tone2<=	7	;
when	139	=>tone2<=	7	;
when	140	=>tone2<=	0	;
when	141	=>tone2<=	8	;
when	142	=>tone2<=	8	;
when	143	=>tone2<=	8	;
when	144	=>tone2<=	8	;
when	145	=>tone2<=	8	;
when	146	=>tone2<=	8	;
when	147	=>tone2<=	0	;
when	148	=>tone2<=	7	;
when	149	=>tone2<=	7	;
when	150	=>tone2<=	0	;
when	151	=>tone2<=	8	;
when	152	=>tone2<=	8	;
when	153	=>tone2<=	8	;
when	154	=>tone2<=	8	;
when	155	=>tone2<=	0	;
when	156	=>tone2<=	10	;
when	157	=>tone2<=	10	;
when	158	=>tone2<=	10	;
when	159	=>tone2<=	10	;
when	160	=>tone2<=	0	;
when	161	=>tone2<=	7	;
when	162	=>tone2<=	7	;
when	163	=>tone2<=	7	;
when	164	=>tone2<=	7	;
when	165	=>tone2<=	7	;
when	166	=>tone2<=	7	;
when	167	=>tone2<=	0	;
when	168	=>tone2<=	3	;
when	169	=>tone2<=	3	;
when	170	=>tone2<=	3	;
when	171	=>tone2<=	3	;
when	172	=>tone2<=	0	;
when	173	=>tone2<=	6	;
when	174	=>tone2<=	6	;
when	175	=>tone2<=	6	;
when	176	=>tone2<=	6	;
when	177	=>tone2<=	6	;
when	178	=>tone2<=	6	;
when	179	=>tone2<=	0	;
when	180	=>tone2<=	5	;
when	181	=>tone2<=	5	;
when	182	=>tone2<=	0	;
when	183	=>tone2<=	6	;
when	184	=>tone2<=	6	;
when	185	=>tone2<=	6	;
when	186	=>tone2<=	6	;
when	187	=>tone2<=	0	;
when	188	=>tone2<=	8	;
when	189	=>tone2<=	8	;
when	190	=>tone2<=	8	;
when	191	=>tone2<=	8	;
when	192	=>tone2<=	0	;
when	193	=>tone2<=	5	;
when	194	=>tone2<=	5	;
when	195	=>tone2<=	5	;
when	196	=>tone2<=	5	;
when	197	=>tone2<=	5	;
when	198	=>tone2<=	5	;
when	199	=>tone2<=	0	;
when	200	=>tone2<=	3	;
when	201	=>tone2<=	3	;
when	202	=>tone2<=	3	;
when	203	=>tone2<=	3	;
when	204	=>tone2<=	0	;
when	205	=>tone2<=	4	;
when	206	=>tone2<=	4	;
when	207	=>tone2<=	4	;
when	208	=>tone2<=	4	;
when	209	=>tone2<=	0	;
when	210	=>tone2<=	8	;
when	211	=>tone2<=	8	;
when	212	=>tone2<=	0	;
when	213	=>tone2<=	7	;
when	214	=>tone2<=	7	;
when	215	=>tone2<=	7	;
when	216	=>tone2<=	7	;
when	217	=>tone2<=	7	;
when	218	=>tone2<=	7	;
when	219	=>tone2<=	0	;
when	220	=>tone2<=	8	;
when	221	=>tone2<=	8	;
when	222	=>tone2<=	8	;
when	223	=>tone2<=	8	;
when	224	=>tone2<=	0	;
when	225	=>tone2<=	9	;
when	226	=>tone2<=	9	;
when	227	=>tone2<=	9	;
when	228	=>tone2<=	9	;
when others =>tone2<=0;
end case;
end case;
end if;
end if;
end process;
end song_arch;